----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:18:21 01/17/2013 
-- Design Name: 
-- Module Name:    main - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SevSegConv is
    Port ( input : in  STD_LOGIC_VECTOR (3 downto 0);
           output : out  STD_LOGIC_VECTOR (6 downto 0)
			  );
end SevSegConv;

architecture Behavioral of SevSegConv is
begin
process(input)
	begin
	case input is
	when  "0000"=> output <= "0000001";
	when  "0001"=> output <= "1001111";
	when  "0010"=> output <= "0010010";
	when  "0011"=> output <= "0000110";
	when  "0100"=> output <= "1001100";
	when  "0101"=> output <= "0100100";
	when  "0110"=> output <= "0100000";
	when  "0111"=> output <= "0001101";
	when  "1000"=> output <= "0000000";
	when  "1001"=> output <= "0000100";
	when  "1010"=> output <= "0001000";
	when  "1011"=> output <= "1100000";
	when  "1100"=> output <= "0110001";
	when  "1101"=> output <= "1000010";
	when  "1110"=> output <= "0110000";
	when  others => output <= "1111111";
	end case;
end process;
end Behavioral;

